// Pipelined Risc-V CPU //
