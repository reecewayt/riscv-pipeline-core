// Testbench for Pipelined Risc-V CPU //

