module decode_unit(

); 
    import riscv_pkg::*;


endmodule: decode_unit